module Loto (Clk, BPBack, BPReview, BPReset, BPTirage, A1, A2, A3, A4); 

input Clk, BPBack, BPReview, BPReset, BPTirage; 

output [6:0] A1; 

output [6:0] A2; 

output [6:0] A3; 

output [6:0] A4; 

 

wire [6:0] A, [6:0] B, [6:0] C, [6:0] D, [6:0] E, [6:0] F, [6:0] G, [6:0] H, [6:0] I, [6:0] J; 

endmodule